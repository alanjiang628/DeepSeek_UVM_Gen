`ifndef __SC_DEFINES_SV__
`define __SC_DEFINES_SV__
`define DEBOUNCE_THRESHOLD 10
`define SRC 3
`endif